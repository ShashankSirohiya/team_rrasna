module axi_lite_read_tb;

endmodule : axi_lite_read_tb